module packet_segmenter #(
  parameter MTU = 64,
  parameter AXI_FRAME_SIZE = 128
  )
  (
  //! INPUTS/OUTPUTS
  input logic clk, rst,
  
  input logic [AXI_FRAME_SIZE-1:0] s_axis_tdata,
  input logic s_axis_tvalid,
  output logic s_axis_tready,
  input logic s_axis_tlast,

  output logic [MTU-1:0] m_axis_tdata,
  output logic m_axis_tvalid,
  input logic m_axis_tready,
  output logic m_axis_tlast
  );

  // HELPER FUNCTIONS

  //Greatest Common Divisor
  function automatic int gcd(input int a, input int b);
    while (b != 0) begin
      int temp = b;
      b = a % b;
      a = temp;
    end
    return a;
  endfunction

  //Lowest Common Multiple
  function automatic int lcm(input int a, input int b);
    if (a == 0 || b == 0)
      return 0;
    else 
      return (a / gcd(a, b)) * b;
  endfunction
  
  initial begin
  assert (AXI_FRAME_SIZE == 128)
    else $warning("Non-standard AXI width for video; 128-bit expected");
  assert (MTU > 0 && MTU <= 128 && (128 % MTU == 0))
    else $warning("MTU should divide 128 for clean video packing");
  end

  generate 
  if (MTU == AXI_FRAME_SIZE) begin : BUFFER_BYPASS
    assign m_axis_tdata = s_axis_tdata;
    assign m_axis_tvalid = s_axis_tvalid;
    assign s_axis_tready = m_axis_tready;
    assign m_axis_tlast = s_axis_tlast;
  end : BUFFER_BYPASS 
  else begin : BUFFER_PATH
    // INTERNAL VARIABLES
    localparam int LCM = lcm(AXI_FRAME_SIZE, MTU);
    logic [LCM-1:0]                        buffer;
    logic [$clog2(LCM/AXI_FRAME_SIZE)-1:0] write_ptr;  
    logic [$clog2(LCM/MTU)-1:0]            read_ptr;
    logic [$clog2(LCM):0]                  bits_stored;

    logic input_last_seen;
    logic [$clog2(LCM/MTU)-1:0] packets_remaining;
            
    // PROCESSES
    always_ff @(posedge clk) begin
      if (rst) begin
        write_ptr <= '0;
        read_ptr <= '0;
        bits_stored <= '0;
        input_last_seen <= '0;
        packets_remaining <= '0;
    end else begin
      if (s_axis_tvalid && s_axis_tready && s_axis_tlast) begin
        input_last_seen <= 1'b1;
        packets_remaining <= ((bits_stored + AXI_FRAME_SIZE) + MTU - 1 ) / MTU;
      end

      if (m_axis_tvalid && m_axis_tready && m_axis_tlast) begin
        input_last_seen <= 1'b0;
        packets_remaining <= '0;
      end

      case ({(m_axis_tvalid), (s_axis_tready && s_axis_tvalid && m_axis_tready)})
      //[1]: read, [0]: write 
        2'b01: begin 
          bits_stored <= bits_stored + AXI_FRAME_SIZE; // write only 
          write_ptr <= (write_ptr >= LCM/AXI_FRAME_SIZE - 1) ? 0 : write_ptr + 1;
        end
        2'b10: begin 
          bits_stored <= bits_stored - MTU; // read only 
          read_ptr <= (read_ptr >= LCM/MTU - 1) ? 0 : read_ptr + 1;
          if (packets_remaining > 0)
            packets_remaining <= packets_remaining - 1;
        end
        2'b11: begin 
          bits_stored <= bits_stored + AXI_FRAME_SIZE - MTU; // read & write
          write_ptr <= (write_ptr >= LCM/AXI_FRAME_SIZE - 1) ? 0 : write_ptr + 1;
          read_ptr <= (read_ptr >= LCM/MTU - 1) ? 0 : read_ptr + 1;
          if (packets_remaining > 0)
            packets_remaining <= packets_remaining - 1;
        end
      endcase

      if (s_axis_tready && s_axis_tvalid && m_axis_tready) begin
        // write to buffer 
        buffer[write_ptr * AXI_FRAME_SIZE +: AXI_FRAME_SIZE] <= s_axis_tdata;
      end
    end

    end

    assign s_axis_tready = (bits_stored + AXI_FRAME_SIZE) <= LCM;
    assign m_axis_tdata = buffer[read_ptr * MTU +: MTU] & {MTU{m_axis_tvalid}};     
    assign m_axis_tvalid = (bits_stored>=MTU) || (input_last_seen && packets_remaining > 0);
    assign m_axis_tlast = input_last_seen && (packets_remaining == 1);

  end : BUFFER_PATH
  endgenerate 
endmodule
